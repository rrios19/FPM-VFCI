// Tecnologico de Costa Rica
// Verificacion funcional de circuitos integrados
// S2 2022
// Proyecto 2: Floating point multipliers
// Irene Prieto 
// Ronald Rios
