// Tecnologico de Costa Rica
// Verificacion funcional de circuitos integrados
// S2 2022
// Project 2: Floating point multipliers
// Irene Prieto 
// Ronald Rios

class example extends uvm_example_something;
	`uvm_object_utils(example); // Register at the factory

	function new(string name = "example"); // Builder
		super.new(name);
	endfunction

	// Your code here
endclass


//:%s/example/newname
